/*
 * Copyright 2023 BSC*
 * *Barcelona Supercomputing Center (BSC)
 * 
 * SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
 * 
 * Licensed under the Solderpad Hardware License v 2.1 (the “License”); you
 * may not use this file except in compliance with the License, or, at your
 * option, the Apache License version 2.0. You may obtain a copy of the
 * License at
 * 
 * https://solderpad.org/licenses/SHL-2.1/
 * 
 * Unless required by applicable law or agreed to in writing, any work
 * distributed under the License is distributed on an “AS IS” BASIS, WITHOUT
 * WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the
 * License for the specific language governing permissions and limitations
 * under the License.
 */

//-----------------------------
// includes
//-----------------------------

`timescale 1 ns / 1 ns
//`default_nettype none

`include "colors.vh"

import drac_pkg::*;

module tb_regfile();

//-----------------------------
// Local parameters
//-----------------------------
    parameter VERBOSE         = 1;
    parameter CLK_PERIOD      = 2;
    parameter CLK_HALF_PERIOD = CLK_PERIOD / 2;

//-----------------------------
// Signals
//-----------------------------
    reg     tb_clk_i;

    logic     [NUM_SCALAR_INSTR-1:0] tb_write_enable_i;
    phreg_t   [NUM_SCALAR_INSTR-1:0] tb_write_addr_i;
    bus64_t [NUM_SCALAR_INSTR-1:0] tb_write_data_i;
    // read ports input
    phreg_t   [NUM_SCALAR_INSTR-1:0] tb_read_addr1_S_i ;
    phreg_t   [NUM_SCALAR_INSTR-1:0] tb_read_addr2_S_i ;
    // read port output
    bus64_t [NUM_SCALAR_INSTR-1:0] tb_read_data1_S_o ;
    bus64_t [NUM_SCALAR_INSTR-1:0] tb_read_data2_S_o ;


//-----------------------------
// Module
//-----------------------------

    regfile regfile_inst( 
        .clk_i(tb_clk_i),
        .write_enable_i(tb_write_enable_i),
        .write_addr_i(tb_write_addr_i),
        .write_data_i(tb_write_data_i),
        .read_addr1_S_i(tb_read_addr1_S_i),
        .read_addr2_S_i(tb_read_addr2_S_i),
        .read_data1_S_o(tb_read_data1_S_o),
        .read_data2_S_o(tb_read_data2_S_o)
    );

//-----------------------------
// DUT
//-----------------------------


//***clk_gen***
// A single clock source is used in this design.
    initial tb_clk_i = 1;
    always #CLK_HALF_PERIOD tb_clk_i = !tb_clk_i;


//***task automatic init_sim***
    task automatic init_sim;
        begin
            $display("*** init_sim");
            tb_clk_i <='{default:1};
            tb_write_enable_i<='{default:0};
            tb_write_addr_i<='{default:0};
            tb_write_data_i<='{default:0};
            tb_read_addr1_S_i<='{default:0};
            tb_read_addr2_S_i<='{default:0};
            
            $display("Done");
            
        end
    endtask

//***task automatic init_dump***
//This task dumps the ALL signals of ALL levels of instance dut_example into the test.vcd file
//If you want a subset to modify the parameters of $dumpvars
    task automatic init_dump;
        begin
            $display("*** init_dump");
            $dumpfile("dump_file.vcd");
            $dumpvars(0,regfile_inst);
        end
    endtask

    task automatic tick();
        begin
            //$display("*** tick");
            #CLK_PERIOD;
        end
    endtask


    task automatic test_sim1;
        output int tmp;
        begin
            //$display("*** tick");
            tmp = 0;
	    #CLK_PERIOD;
            tb_write_enable_i = '{NUM_SCALAR_INSTR{1'b1}};
            tb_write_addr_i[0] = 5'b00001;
             tb_write_addr_i[1] = 5'b00010;
            tb_write_data_i = '{NUM_SCALAR_INSTR{64'h01}};
            tb_read_addr1_S_i = '{NUM_SCALAR_INSTR{5'b00000}};
            tb_read_addr2_S_i = '{NUM_SCALAR_INSTR{5'b00000}};
            #CLK_PERIOD;
            tb_write_enable_i = '{NUM_SCALAR_INSTR{1'b0}};
	        tb_write_addr_i = '{NUM_SCALAR_INSTR{5'b00000}};
            for(int i=0;i<NUM_SCALAR_INSTR;i++) begin
            assert(tb_read_data1_S_o[i] == 0) else begin tmp++; assert(1 == 0); end
            assert(tb_read_data2_S_o[i] == 0) else begin tmp++; assert(1 == 0); end
            tb_read_addr1_S_i[i] = 5'b00001;
            tb_read_addr2_S_i[i] = 5'b00001;
            end
	    #CLK_PERIOD;
         for(int i=0;i<NUM_SCALAR_INSTR;i++) begin
            assert(tb_read_data1_S_o[i] == 64'h01) else begin tmp++; assert(1 == 0); end
            assert(tb_read_data2_S_o[i] == 64'h01) else begin tmp++; assert(1 == 0); end
         end
        end
    endtask

//***task automatic test_sim***
    task automatic test_sim;
        begin
            int tmp;
            $display("*** test_sim");
            test_sim1(tmp);
	    if(tmp == 0) begin
                `START_GREEN_PRINT
                $display("PASS");
                `END_COLOR_PRINT
	    end else begin
                `START_RED_PRINT
                $error("FAIL");
                `END_COLOR_PRINT
            end
        end
    endtask


//***init_sim***
//The tasks that compose my testbench are executed here, feel free to add more tasks.
    initial begin
        init_sim();
        init_dump();
        test_sim();
    end


endmodule
//`default_nettype wire
